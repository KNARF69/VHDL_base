library ieee;
use ieee.std_logic_1164.all;

entity fpga_io_tort is
    generic (

        
    )
